`define RB 2'b00
`define RADD 2'b01
`define RSUB 2'b10
`define RMULT 2'b11