`define NOP 3'b010
`define ADD 3'b001
`define MULT 3'b011
`define ADDI 3'b101
`define COPY 3'b110
`define MULTI 3'b111
`define WLD0 3'b000 // Wait for SW9=0 then load into register
`define WLD1 3'b100 // Wait for SW9=1 then load into register