`define DATA_BUS_SIZE 8
`define INSTRUCTION_SIZE 14
`define PROGRAM_CODE_SIZE 4 // up to 16 instructions
`define REGISTERS_SIZE 3 // 8 registers
`define ALU_CODE_SIZE 2 // up to 4 alu codes
`define OPCODE_SIZE 3 // up to 8 opcodes